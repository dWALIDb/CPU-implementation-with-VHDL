library IEEE;
use ieee.std_logic_1164.all;
use work.tools.all;

entity cu is 
port 
(
	--status of our micro processor
	flag_reg:in std_logic_vector(dataBus_size-1 downto 0);
	ir_output :in std_logic_vector(dataBus_size-1 downto 0);
	--usual controlers of cu
	clk,reset,int,go:in std_logic;
	-- data path's controlable signals
	RF_address: out	std_logic_vector(RF_adress-1 downto 0);
	alu_op: 	out std_logic_vector(alu_ops-1 downto 0);
	shifter_op: out std_logic_vector(shifter_ops-1 downto 0);
	to_freg : 	out std_logic_vector(0 downto 0);
	to_acc_sel,to_RF_sel,memory_data_sel: out std_logic_vector(1 downto 0);
	carry_sel,rf_read,rf_write: out std_logic;
	acc_enable,freg_enable,swap_reg_enable: out std_logic;
	-- memory's controlable signals
	spc_sel:out std_logic_vector(0 downto 0);
	ir_adress:out std_logic_vector(1 downto 0);
	pc_enable,ix_enable,mar_enable,mir_enable,sp_enable,ram_enable: out std_logic;
	au_op:out std_logic_vector(1 downto 0);
	au_in_sel,mir_sel,mar_sel:out std_logic_vector(1 downto 0);
	ram_read,ram_write,ir_read,ir_write: out std_logic;
	-- io port's controlable signals 
	io_sel: out std_logic_vector(0 downto 0);
	io_wd,io_rd,io_write: out std_logic;
	io_adress:out std_logic_vector(3 downto 0)
);
end cu;
architecture arch of cu is

signal microinstruction: opcodes:=fetch;
signal current_instruction: std_logic_vector(dataBus_size-1 downto 0);
signal int_enable:std_logic:='0';
signal t_state:integer range 0 to 12;
signal go_next:boolean:=false;
signal control:std_logic_vector(49 downto 0);

begin
next_state:	process(clk,reset,int_enable,go_next,go)
	begin
	if reset='1' then microinstruction<=fetch;
	elsif (clk'event and clk='0' and go_next=true and go='1') then 
	case microinstruction is 
	when fetch=> current_instruction<=ir_output;--we need to keep opcode since ir changes and sends different data to cu
	microinstruction<=decode;
	when decode=>
		case(current_instruction)is 
		when x"00"=>microinstruction<=ldd  ;when x"17"=>microinstruction<=rotr ;when x"2E"=>microinstruction<=jr    ;	when x"46"=>microinstruction<=jpn	  ;when x"5D"=>microinstruction<=incrc;
		when x"01"=>microinstruction<=ldr  ;when x"18"=>microinstruction<=adr  ;when x"2F"=>microinstruction<=jpe   ;	when x"47"=>microinstruction<=jpo 	  ;when x"5E"=>microinstruction<=decrc;
		when x"02"=>microinstruction<=ldi  ;when x"19"=>microinstruction<=adm  ;when x"30"=>microinstruction<=jpl   ;	when x"48"=>microinstruction<=jpno 	  ;when x"5F"=>microinstruction<=incz;
		when x"03"=>microinstruction<=rla  ;when x"1A"=>microinstruction<=adi  ;when x"31"=>microinstruction<=jpg   ;	when x"49"=>microinstruction<=jrc 	  ;when x"60"=>microinstruction<=decz;
											when x"1B"=>microinstruction<=sbr  ;when x"32"=>microinstruction<=jre   ;	when x"4A"=>microinstruction<=jrnc 	  ;when x"61"=>microinstruction<=incrz;
		when x"05"=>microinstruction<=rli  ;when x"1C"=>microinstruction<=sbm  ;when x"33"=>microinstruction<=jrl   ;	when x"4B"=>microinstruction<=jrz	  ;when x"62"=>microinstruction<=decrz;
		when x"06"=>microinstruction<=rlm  ;when x"1D"=>microinstruction<=sbi  ;when x"34"=>microinstruction<=jrg   ;	when x"4C"=>microinstruction<=jrnz 	  ;when x"63"=>microinstruction<=adix;
		when x"07"=>microinstruction<=sta  ;when x"1E"=>microinstruction<=swp  ;when x"35"=>microinstruction<=jpne  ;	when x"4D"=>microinstruction<=jrp 	  ;when x"64"=>microinstruction<=sbix;
		when x"08"=>microinstruction<=str  										;when x"36"=>microinstruction<=jrne  ;when x"4E"=>microinstruction<=jrn 	  ;when x"65"=>microinstruction<=andix;
		when x"09"=>microinstruction<=ldsp ;when x"20"=>microinstruction<=incix ;when x"37"=>microinstruction<=jpc   ;	when x"4F"=>microinstruction<=jro 	  ;when x"66"=>microinstruction<=orix;
		when x"0A"=>microinstruction<=ldix ;when x"21"=>microinstruction<=decix ;when x"38"=>microinstruction<=jpnc  ;	when x"50"=>microinstruction<=jrno 	  ;when x"67"=>microinstruction<=xorix;
		when x"0B"=>microinstruction<=inc  ;when x"22"=>microinstruction<=andr ;when x"39"=>microinstruction<=jpz   ;	when x"51"=>microinstruction<=pushacc ;when x"68"=>microinstruction<=cpix;
		when x"0C"=>microinstruction<=incr ;when x"23"=>microinstruction<=andm ;when x"3A"=>microinstruction<=jpnz  ;	when x"52"=>microinstruction<=popacc  ;when x"69"=>microinstruction<=pctoix;
		when x"0D"=>microinstruction<=dec  ;when x"24"=>microinstruction<=andi ;when x"3B"=>microinstruction<=jpp   ;	when x"53"=>microinstruction<=pushreg ;when x"6A"=>microinstruction<=offsetix;
		when x"0E"=>microinstruction<=decr ;when x"25"=>microinstruction<=orr  ;when x"3C"=>microinstruction<=call  ;	when x"54"=>microinstruction<=popreg  ;when x"6B"=>microinstruction<=pushix;
		when x"0F"=>microinstruction<=cp   ;when x"26"=>microinstruction<=orm  ;when x"55"=>microinstruction<=di    ;   when x"3E"=>microinstruction<=ret;     when x"6C"=>microinstruction<=popix;
		when x"10"=>microinstruction<=cpr  ;when x"27"=>microinstruction<=ori  ;when x"56"=>microinstruction<=ei	 ;  when x"3F"=>microinstruction<=pushflag;
		when x"11"=>microinstruction<=cpm  ;when x"28"=>microinstruction<=xorr ;when x"57"=>microinstruction<=ina     ; when x"40"=>microinstruction<=popflag; 
		when x"12"=>microinstruction<=sl   ;when x"29"=>microinstruction<=xorm ;when x"58"=>microinstruction<=inr 	  ; when x"41"=>microinstruction<=indexedld;
		when x"13"=>microinstruction<=sr   ;when x"2A"=>microinstruction<=xori ;when x"59"=>microinstruction<=outa 	  ; when x"42"=>microinstruction<=indexedstr;
		when x"14"=>microinstruction<=rot  ;when x"2B"=>microinstruction<=cpl  ;when x"5A"=>microinstruction<=outr 	  ; when x"43"=>microinstruction<=get;
		when x"15"=>microinstruction<=slr  ;when x"2C"=>microinstruction<=neg  ;when x"FF"=>microinstruction<=halt ;    when x"5B"=>microinstruction<=incc;
		when x"16"=>microinstruction<=srr  ;when x"2D"=>microinstruction<=jp   ;when x"5C"=>microinstruction<=decc;	when OTHERS=>microinstruction<=nop ;
			end case;
	when ldd  => nextstate(int,int_enable,microinstruction);when rotr => nextstate(int,int_enable,microinstruction);when jpn	 => nextstate(int,int_enable,microinstruction);when jr    => nextstate(int,int_enable,microinstruction);when decc=>nextstate(int,int_enable,microinstruction);
	when ldr  => nextstate(int,int_enable,microinstruction);when adr  => nextstate(int,int_enable,microinstruction);when jpo 	 => nextstate(int,int_enable,microinstruction);when jpe   => nextstate(int,int_enable,microinstruction);when incrc=>nextstate(int,int_enable,microinstruction);
	when ldi  => nextstate(int,int_enable,microinstruction);when adm  => nextstate(int,int_enable,microinstruction);when jpno 	 => nextstate(int,int_enable,microinstruction);when jpl   => nextstate(int,int_enable,microinstruction);when decrc=>nextstate(int,int_enable,microinstruction);
	when rla  => nextstate(int,int_enable,microinstruction);when adi  => nextstate(int,int_enable,microinstruction);when jrc 	 => nextstate(int,int_enable,microinstruction);when jpg   => nextstate(int,int_enable,microinstruction);when incz=>nextstate(int,int_enable,microinstruction);
	when sbr  => nextstate(int,int_enable,microinstruction);when jrnc 	 => nextstate(int,int_enable,microinstruction);when jre   => nextstate(int,int_enable,microinstruction);
	when rli  => nextstate(int,int_enable,microinstruction);when sbm  => nextstate(int,int_enable,microinstruction);when jrz	 => nextstate(int,int_enable,microinstruction);when jrl   => nextstate(int,int_enable,microinstruction);when decz=>nextstate(int,int_enable,microinstruction);
	when rlm  => nextstate(int,int_enable,microinstruction);when sbi  => nextstate(int,int_enable,microinstruction);when jrnz 	 => nextstate(int,int_enable,microinstruction);when jrg   => nextstate(int,int_enable,microinstruction);when incrz=>nextstate(int,int_enable,microinstruction);
	when sta  => nextstate(int,int_enable,microinstruction);when swp  => nextstate(int,int_enable,microinstruction);when jrp 	 => nextstate(int,int_enable,microinstruction);when jpne  => nextstate(int,int_enable,microinstruction);when decrz=>nextstate(int,int_enable,microinstruction);
	when str  => nextstate(int,int_enable,microinstruction);when nop  => nextstate(int,int_enable,microinstruction);when jrn 	 => nextstate(int,int_enable,microinstruction);when jrne  => nextstate(int,int_enable,microinstruction);when adix=>nextstate(int,int_enable,microinstruction);
	when ldsp => nextstate(int,int_enable,microinstruction);when incix=> nextstate(int,int_enable,microinstruction);when jro 	 => nextstate(int,int_enable,microinstruction);when jpc   => nextstate(int,int_enable,microinstruction);when sbix=>nextstate(int,int_enable,microinstruction);
	when ldix => nextstate(int,int_enable,microinstruction);when decix=> nextstate(int,int_enable,microinstruction);when jrno 	 => nextstate(int,int_enable,microinstruction);when jpnc  => nextstate(int,int_enable,microinstruction);when orix=>nextstate(int,int_enable,microinstruction);
	when inc  => nextstate(int,int_enable,microinstruction);when andr => nextstate(int,int_enable,microinstruction);when pushacc => nextstate(int,int_enable,microinstruction);when jpz   => nextstate(int,int_enable,microinstruction);when andix=>nextstate(int,int_enable,microinstruction);
	when incr => nextstate(int,int_enable,microinstruction);when andm => nextstate(int,int_enable,microinstruction);when popacc  => nextstate(int,int_enable,microinstruction);when jpnz  => nextstate(int,int_enable,microinstruction);when xorix=>nextstate(int,int_enable,microinstruction);
	when dec  => nextstate(int,int_enable,microinstruction);when andi => nextstate(int,int_enable,microinstruction);when pushreg => nextstate(int,int_enable,microinstruction);when jpp   => nextstate(int,int_enable,microinstruction);when cpix=>nextstate(int,int_enable,microinstruction);
	when decr => nextstate(int,int_enable,microinstruction);when orr  => nextstate(int,int_enable,microinstruction);when popreg  => nextstate(int,int_enable,microinstruction);when interrupt=>microinstruction<=fetch;					when pctoix=>nextstate(int,int_enable,microinstruction);
	when cp   => nextstate(int,int_enable,microinstruction);when ori  => nextstate(int,int_enable,microinstruction);when di  	 => nextstate(int,int_enable,microinstruction);when popflag=>nextstate(int,int_enable,microinstruction);when offsetix=>nextstate(int,int_enable,microinstruction);
	when cpr  => nextstate(int,int_enable,microinstruction);when orm  => nextstate(int,int_enable,microinstruction);when ei 	 => nextstate(int,int_enable,microinstruction);when pushflag=>nextstate(int,int_enable,microinstruction);when pushix=>nextstate(int,int_enable,microinstruction);
	when cpm  => nextstate(int,int_enable,microinstruction);when xori => nextstate(int,int_enable,microinstruction);when ina     => nextstate(int,int_enable,microinstruction);when indexedld=>nextstate(int,int_enable,microinstruction);when popix=>nextstate(int,int_enable,microinstruction);
	when sl   => nextstate(int,int_enable,microinstruction);when xorr => nextstate(int,int_enable,microinstruction);when inr 	 => nextstate(int,int_enable,microinstruction);when indexedstr=>nextstate(int,int_enable,microinstruction);
	when sr   => nextstate(int,int_enable,microinstruction);when xorm => nextstate(int,int_enable,microinstruction);when outa 	 => nextstate(int,int_enable,microinstruction);when get=>nextstate(int,int_enable,microinstruction);
	when rot  => nextstate(int,int_enable,microinstruction);when cpl  => nextstate(int,int_enable,microinstruction);when outr 	 => nextstate(int,int_enable,microinstruction);when incc=>nextstate(int,int_enable,microinstruction);
	when slr  => nextstate(int,int_enable,microinstruction);when neg  => nextstate(int,int_enable,microinstruction);when halt 	 => microinstruction<=halt;when call=>nextstate(int,int_enable,microinstruction);when ret=>nextstate(int,int_enable,microinstruction);                 
	when srr  => nextstate(int,int_enable,microinstruction);when jp   => nextstate(int,int_enable,microinstruction);when others=>microinstruction<=nop;
	end case;
	end if;
	end process;
	
output_logic:process(microinstruction,t_state,clk,reset,go,go_next,ir_output,control,flag_reg)
	begin
			--a counter for the T states :)
		if reset='1'or microinstruction=halt  then t_state<=0;
	elsif(clk'event and clk='0' and go='1') then 
		if(go_next=true)then t_state<=0;
			else t_state<=t_state+1; end if;end if;
		
		--set initial conditions for control bus inside CU ;)
		go_next<=false; 

		io_write<='0';

		control<=(others=>'0');

		if (rising_edge(clk) and microinstruction=ei) then int_enable<='1';end if; 
		if(rising_edge(clk) and (microinstruction=interrupt or microinstruction=di)) then int_enable<='0';
		end if;
		--the acctual combinational logic output
	case(microinstruction)is
	when fetch=>if(t_state=0) then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			 elsif(t_state=1) then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			 elsif(t_state=2) then control<="0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
								   go_next<=true; end if;
	when decode=>control<=(others=>'0');go_next<=true;
	when ldd=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"01"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"11"&"0");
			elsif(t_state=3)then control<=("1"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"01"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			go_next<=true;end if;
	when ldr=>if(t_state=0) then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"01"&"00"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"01"&"00"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when ldi=>if(t_state=0) then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"01"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
								   go_next<=true; end if;
	when rla=>if(t_state=0)then  control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"0"&"1"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"01"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
								   go_next<=true;end if;
	when rli=>if(t_state=0) then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=3)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"0"&"1"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
								  go_next<=true;end if;
	when rlm=>if(t_state=0) then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0"); 
			elsif(t_state=3)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"10"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=4)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"10"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"11"&"0");
			elsif(t_state=5)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"0"&"1"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when sta=>if(t_state=0) then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"10"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"1"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"10"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"01"&"11"&"0");
			elsif(t_state=3)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"0"&"1"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when str=>if(t_state=0) then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=3)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"10"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=4)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"10"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"11"&"0");
			elsif(t_state=5)then control<=("0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=6)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"0"&"1"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when ldsp=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when ldix=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when inc=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
		elsif(t_state=1)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0011"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when incc=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
		elsif(t_state=1)then control<=("0"&flag_reg(2)&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0011"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when incz=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
		elsif(t_state=1)then control<=("0"&flag_reg(3)&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0011"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when incr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"1"&"0000"&"0"&"0"&"0100"&"10"&"00"&"0"&"00"&"01"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when incrc=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&flag_reg(2)&"0000"&"0"&"0"&"0100"&"10"&"00"&"0"&"00"&"01"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when incrz=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&flag_reg(3)&"0000"&"0"&"0"&"0100"&"10"&"00"&"0"&"00"&"01"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when dec=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
		elsif(t_state=1)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0101"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when decc=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
		elsif(t_state=1)then control<=("0"&flag_reg(2)&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0101"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when decz=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
		elsif(t_state=1)then control<=("0"&flag_reg(3)&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0101"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when decr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"1"&"0000"&"0"&"0"&"0110"&"10"&"00"&"0"&"00"&"01"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when decrc=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&flag_reg(2)&"0000"&"0"&"0"&"0110"&"10"&"00"&"0"&"00"&"01"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when decrz=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&flag_reg(3)&"0000"&"0"&"0"&"0110"&"10"&"00"&"0"&"00"&"01"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when cp =>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when cpr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when cpm=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"11"&"0");
			elsif(t_state=3)then control<=("1"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when sl=>if(t_state=0) then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"10"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when sr=>if(t_state=0) then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"01"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when rot=>if(t_state=0)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"11"&"0"&"00"&"00"&"00"&"1"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when slr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"1"&"0000"&"0"&"0"&"1100"&"10"&"10"&"0"&"00"&"01"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when srr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"1"&"0000"&"0"&"0"&"1100"&"10"&"01"&"0"&"00"&"01"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when rotr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"1"&"0000"&"0"&"0"&"1100"&"10"&"11"&"0"&"00"&"01"&"10"&"1"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when adr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"0"&"0000"&"0"&"0"&"0001"&"00"&"00"&"0"&"00"&"00"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when adm=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"11"&"0");
			elsif(t_state=3)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0001"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when adi=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0001"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when sbr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"0"&"0000"&"0"&"0"&"0010"&"00"&"00"&"0"&"00"&"00"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when sbm=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"11"&"0");
			elsif(t_state=3)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0010"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when sbi=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0010"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when swp=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=3)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(dataBus_size-2 downto dataBus_size-4)&"0"&"1"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"11"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when incix=>if(t_state=0)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"10"&"00"&"00"&"0");
									go_next<=true;end if;
	when decix=>if(t_state=0)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"11"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"10"&"00"&"00"&"0");
									go_next<=true;end if;
	when andr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"0"&"0000"&"0"&"0"&"0111"&"00"&"00"&"0"&"00"&"00"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when andm=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"11"&"0");
			elsif(t_state=3)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0111"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when andi=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0111"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when orr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"0"&"0000"&"0"&"0"&"1000"&"00"&"00"&"0"&"00"&"00"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when orm=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"11"&"0");
			elsif(t_state=3)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"1000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when ori=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"1000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when xorr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"0"&"0000"&"0"&"0"&"1011"&"00"&"00"&"0"&"00"&"00"&"10"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when xorm=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"11"&"0");
			elsif(t_state=3)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"1011"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when xori=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"1011"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when cpl=>if(t_state=0)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"1001"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when neg=>if(t_state=0)then control<=("0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"1010"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jp=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jpe=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(5)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jpl=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(4)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jpg=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(6)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jpne=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(not flag_reg(5)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jre=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(5)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jrl=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(4)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jrg=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(6)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jrne=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(not flag_reg(5)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jpc=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(2)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jpnc=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(not flag_reg(2)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jpz=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(3)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jpnz=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(not flag_reg(3)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jpp=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(0)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jpn=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(not flag_reg(0)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jpo=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(1)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jpno=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(not flag_reg(1)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jrc=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(2)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jrnc=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(not flag_reg(2)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jrz=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(3)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jrnz=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(not flag_reg(3)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jrp=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(0)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jrn=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(not flag_reg(0)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jro=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(flag_reg(1)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when jrno=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=(not flag_reg(1)&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when pushacc=>if(t_state=0)then control<=("0"&"0"&"1"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"01"&"10"&"0");
				elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"1"&"0"&"1"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"11"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"01"&"00"&"00"&"0");
									go_next<=true;end if;
	when popacc=>if(t_state=0)then control<=("0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"01"&"00"&"00"&"0");
				elsif(t_state=1)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"10"&"0");
				elsif(t_state=2)then control<=("0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"01"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when pushreg=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
				elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
				elsif(t_state=2)then control<=("0"&"0"&"1"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"10"&"0");
				elsif(t_state=3)then control<=("0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"1"&"0"&"1"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"11"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"01"&"00"&"00"&"0");
									go_next<=true;end if;
	when popreg=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"01"&"00"&"00"&"0");
				elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
				elsif(t_state=2)then control<=("1"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"10"&"0");
				elsif(t_state=3)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"0"&"1"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when call=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"1"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"10"&"10"&"0");
			elsif(t_state=3)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"0"&"1"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
			elsif(t_state=4)then control<=("0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"11"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"01"&"00"&"00"&"0");
									go_next<=true;end if;
	when ret=>if(t_state=0)then control<=("0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"01"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"10"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=3)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when di=>if(t_state=0)then go_next<=true;end if;
	when ei=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"11"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
								go_next<=true;end if;
	when ina=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&ir_output(3 downto 0)&"1"&"0"&"0000"&"00"&"00"&"0"&"10"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when outa=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&ir_output(3 downto 0)&"0"&"1"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"1");
									go_next<=true;end if;
	when inr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"0"&"1"&ir_output(dataBus_size-1 downto dataBus_size-4)&"1"&"0"&"0000"&"00"&"00"&"0"&"00"&"10"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when outr=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&ir_output(2 downto 0)&"1"&"0"&ir_output(dataBus_size-1 downto dataBus_size-4)&"0"&"1"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when nop=> control<=(others=>'0');go_next<=true;
	when halt=> control<=(others=>'0');
	when interrupt=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
			elsif(t_state=2)then control<=("0"&"0"&"1"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"10"&"10"&"0");
			elsif(t_state=3)then control<=("1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"0"&"1"&"11"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0");
			elsif(t_state=4)then control<=("0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"11"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"01"&"00"&"00"&"0");
									go_next<=true;end if;
	when pushflag=>if(t_state=0)then control<=("0"&"0"&"1"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"11"&"10"&"0");
				elsif(t_state=1)then control<=("0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"1"&"0"&"1"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"11"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"01"&"00"&"00"&"0");
									go_next<=true;end if;
	when popflag=>if(t_state=0)then control<=("0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"01"&"00"&"10"&"0");
				elsif(t_state=1)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"10"&"0");
				elsif(t_state=2)then control<=("0"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"1"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when indexedld=>if(t_state=0)then control<=("0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"01"&"0");
				elsif(t_state=1)then  control<=("0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"01"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0");
									go_next<=true;end if;
	when indexedstr=>if(t_state=0)then control<=("0"&"0"&"1"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"01"&"01"&"0");
				elsif(t_state=1)then   control<=("0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"0"&"1"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0"); 
									go_next<=true;end if;
	when get=>io_write<='1';if(t_state=0)then control<="0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
			elsif(t_state=1)then control<="1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
			elsif(t_state=2)then control<="0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&ir_output(3 downto 0)&"0"&"1"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"01"&"0";
									go_next<=true;end if;
	when adix=>if(t_state=0)then control<="0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"01"&"0";
			elsif(t_state=1)then control<="0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0001"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
									go_next<=true;end if;
	when sbix=>if(t_state=0)then control<="0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"01"&"0";
			elsif(t_state=1)then control<="0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0010"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
									go_next<=true;end if;
	when andix=>if(t_state=0)then control<="0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"01"&"0";
			elsif(t_state=1)then control<="0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0111"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
									go_next<=true;end if;
	when orix=>if(t_state=0)then control<="0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"01"&"0";
			elsif(t_state=1)then control<="0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"1000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
									go_next<=true;end if;
	when xorix=>if(t_state=0)then control<="0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"01"&"0";
			elsif(t_state=1)then control<="0"&"1"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"1011"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
									go_next<=true;end if;
	when cpix=>if(t_state=0)then control<="0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"01"&"0";
			 elsif(t_state=1)then control<="0"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"01"&"0";
									go_next<=true;end if;
	when pctoix=>if(t_state=0)then control<="0"&"0"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
									go_next<=true;end if;
	when offsetix=>if(t_state=0)then control<="0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
				 elsif(t_state=1)then control<="1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"00"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
				 elsif(t_state=2)then control<="0"&"0"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"00"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"01"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"10"&"00"&"00"&"0";
									go_next<=true;end if;
	when pushix=>if(t_state=0)then control<="0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"11"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"01"&"00"&"00"&"0";
			  elsif(t_state=1)then control<="0"&"0"&"1"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"10"&"10"&"0";
			  elsif(t_state=2)then control<="0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"1"&"0"&"1"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"01"&"00"&"00"&"0";
			  elsif(t_state=3)then control<="1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"10"&"00"&"00"&"0";
			  elsif(t_state=4)then control<="0"&"0"&"1"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"10"&"10"&"0";
			  elsif(t_state=5)then control<="0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"1"&"0"&"1"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"11"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"01"&"00"&"00"&"0";
			  elsif(t_state=6)then control<="0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"10"&"0";
			  elsif(t_state=7)then control<="0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
			  elsif(t_state=8)then control<="1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0";
									go_next<=true;end if;
	when popix=>if(t_state=0) then control<="0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"10"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"01"&"00"&"00"&"0";
			  elsif(t_state=1)then control<="0"&"0"&"1"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"10"&"0";
			  elsif(t_state=2)then control<="0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"0"&"1"&"00"&"0"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
			  elsif(t_state=3)then control<="0"&"0"&"0"&"0"&"0"&"0"&"0"&"0"&"1"&"1"&"0"&"01"&"0"&"1"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"0"&"00"&"00"&"00"&"0";
			  elsif(t_state=4)then control<="0"&"0"&"0"&"0"&"0"&"0"&"1"&"0"&"0"&"0"&"0"&"01"&"1"&"0"&"000"&"0"&"0"&"0000"&"0"&"0"&"0000"&"00"&"00"&"0"&"00"&"00"&"00"&"0"&"1"&"00"&"00"&"00"&"0";
									go_next<=true;end if;
	when others=>control<=(others=>'0');
	end case;

	end process;
	state_out(control,RF_address,alu_op,shifter_op,to_freg,to_acc_sel,to_RF_sel,memory_data_sel,carry_sel,rf_read,rf_write,acc_enable,freg_enable,swap_reg_enable,spc_sel,ir_adress,pc_enable,ix_enable,
	mar_enable,mir_enable,sp_enable,ram_enable,au_op,au_in_sel,mir_sel,mar_sel,ram_read,ram_write,ir_read,ir_write,io_sel,io_wd,io_rd,io_adress);
	

end arch;

